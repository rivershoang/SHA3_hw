import keccak_pkg::plane;
import keccak_pkg::state;
import keccak_pkg::N;

module array_to_string (
	input  state A ,
	output logic [1599:0] S
);
   always_comb begin
   S[63:0] 	= A[0][0];
   S[127:64] 	= A[0][1]; 
   S[191:128]	= A[0][2];
   S[255:192]	= A[0][3];
   S[319:256]	= A[0][4];

   S[383:320]	= A[1][0];
   S[447:384]	= A[1][1];
   S[511:448]	= A[1][2];
   S[575:512]	= A[1][3];
   S[639:576]	= A[1][4];

   S[703:640]	= A[2][0];
   S[767:704]	= A[2][1];
   S[831:768]	= A[2][2];
   S[895:832]	= A[2][3];
   S[959:896]	= A[2][4];

   S[1023:960]	= A[3][0];
   S[1087:1024]	= A[3][1];
   S[1151:1088]	= A[3][2];
   S[1215:1152]	= A[3][3];
   S[1279:1216]	= A[3][4];

   S[1343:1280]	= A[4][0];
   S[1407:1344]	= A[4][1];
   S[1471:1408]	= A[4][2];
   S[1535:1472]	= A[4][3];
   S[1599:1536]	= A[4][4];
   end

endmodule